`timescale 1ns / 1ps
module And(
	input in1,
	input in2,
	output out
   );
	assign out=in1&in2;
endmodule
